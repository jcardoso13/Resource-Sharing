library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity control_unit is

port(
	clk: in std_logic;
	rst: in std_logic
);

end control_unit;


architecture Behavioral of control_unit is


end Behavioral;
